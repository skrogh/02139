library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
entity rom is
port( addr : in std_logic_vector( 9 downto 0 );
do : out std_logic_vector( 12 downto 0 ) );
end rom;
architecture behavioural of rom is
begin
with addr select
do <= "1101111100100" WHEN "0000000000",
"0011001100100" WHEN "0000000001",
"1001001101001" WHEN "0000000010",
"0010110110001" WHEN "0000000011",
"0110010000101" WHEN "0000000100",
"0101110010001" WHEN "0000000101",
"0110100110000" WHEN "0000000110",
"1001111001101" WHEN "0000000111",
"0000001111110" WHEN "0000001000",
"0101111001110" WHEN "0000001001",
"0100110010011" WHEN "0000001010",
"0000001101011" WHEN "0000001011",
"0011010111101" WHEN "0000001100",
"0001110100111" WHEN "0000001101",
"0111110100110" WHEN "0000001110",
"0101000011101" WHEN "0000001111",
"0011001100001" WHEN "0000010000",
"0000101100000" WHEN "0000010001",
"1001000100111" WHEN "0000010010",
"0110010000011" WHEN "0000010011",
"0111100110001" WHEN "0000010100",
"1001001000111" WHEN "0000010101",
"1111101011000" WHEN "0000010110",
"1111001000000" WHEN "0000010111",
"1100110110000" WHEN "0000011000",
"0110011000101" WHEN "0000011001",
"1100111110110" WHEN "0000011010",
"0011000100110" WHEN "0000011011",
"0001100010111" WHEN "0000011100",
"1101101011011" WHEN "0000011101",
"1000101101001" WHEN "0000011110",
"0101101011100" WHEN "0000011111",
"1000110001100" WHEN "0000100000",
"0000000001010" WHEN "0000100001",
"0100011111110" WHEN "0000100010",
"0010000001010" WHEN "0000100011",
"0011000000110" WHEN "0000100100",
"1110000001010" WHEN "0000100101",
"1111101100101" WHEN "0000100110",
"1011011001001" WHEN "0000100111",
"1001100111010" WHEN "0000101000",
"1110011001001" WHEN "0000101001",
"1001001000100" WHEN "0000101010",
"0010100001111" WHEN "0000101011",
"1110000001000" WHEN "0000101100",
"0010110100000" WHEN "0000101101",
"0110101000000" WHEN "0000101110",
"0011101010100" WHEN "0000101111",
"1111111101001" WHEN "0000110000",
"0010011100010" WHEN "0000110001",
"1000001000110" WHEN "0000110010",
"0011110110010" WHEN "0000110011",
"1100011010101" WHEN "0000110100",
"1101100011110" WHEN "0000110101",
"1111010001101" WHEN "0000110110",
"1110001101000" WHEN "0000110111",
"0010000110001" WHEN "0000111000",
"1010011100110" WHEN "0000111001",
"1011000111000" WHEN "0000111010",
"0100101110000" WHEN "0000111011",
"1111101011100" WHEN "0000111100",
"1000101111110" WHEN "0000111101",
"0100000000100" WHEN "0000111110",
"0011100111010" WHEN "0000111111",
"0100001100111" WHEN "0001000000",
"0110001000101" WHEN "0001000001",
"0011100011011" WHEN "0001000010",
"1010001000001" WHEN "0001000011",
"1010010101110" WHEN "0001000100",
"1101011011110" WHEN "0001000101",
"1001001110001" WHEN "0001000110",
"1000000011001" WHEN "0001000111",
"0100011101001" WHEN "0001001000",
"0111101110000" WHEN "0001001001",
"0101111010101" WHEN "0001001010",
"0100001001000" WHEN "0001001011",
"1000101110101" WHEN "0001001100",
"0110010011100" WHEN "0001001101",
"0110000111101" WHEN "0001001110",
"1101000000111" WHEN "0001001111",
"0010110000111" WHEN "0001010000",
"1100000000011" WHEN "0001010001",
"0100101101100" WHEN "0001010010",
"1011111011011" WHEN "0001010011",
"0010100010001" WHEN "0001010100",
"1100010010110" WHEN "0001010101",
"0111010100011" WHEN "0001010110",
"1111010101111" WHEN "0001010111",
"1111100100000" WHEN "0001011000",
"0111100011100" WHEN "0001011001",
"0000001111101" WHEN "0001011010",
"1001111110010" WHEN "0001011011",
"0010110000010" WHEN "0001011100",
"1100110100110" WHEN "0001011101",
"0001110110110" WHEN "0001011110",
"0010011100110" WHEN "0001011111",
"0001010011010" WHEN "0001100000",
"1011000000100" WHEN "0001100001",
"0011100011001" WHEN "0001100010",
"0111100111101" WHEN "0001100011",
"0111100110101" WHEN "0001100100",
"1101101110101" WHEN "0001100101",
"0001001011001" WHEN "0001100110",
"1101111001011" WHEN "0001100111",
"0100001010100" WHEN "0001101000",
"0100100111011" WHEN "0001101001",
"1011000100010" WHEN "0001101010",
"0010111100000" WHEN "0001101011",
"1111111011100" WHEN "0001101100",
"0110111010011" WHEN "0001101101",
"1110101000100" WHEN "0001101110",
"0110010110011" WHEN "0001101111",
"1011100101000" WHEN "0001110000",
"1001000011000" WHEN "0001110001",
"0101101000001" WHEN "0001110010",
"0000000001000" WHEN "0001110011",
"1111101110011" WHEN "0001110100",
"1101110100001" WHEN "0001110101",
"0101000111100" WHEN "0001110110",
"1110111110010" WHEN "0001110111",
"0001000110101" WHEN "0001111000",
"0001100010110" WHEN "0001111001",
"0100010100101" WHEN "0001111010",
"0110101111100" WHEN "0001111011",
"1001010000000" WHEN "0001111100",
"0010110000100" WHEN "0001111101",
"0111010011111" WHEN "0001111110",
"0100010101100" WHEN "0001111111",
"0000001101111" WHEN "0010000000",
"0001011100100" WHEN "0010000001",
"0001110100000" WHEN "0010000010",
"0000000110010" WHEN "0010000011",
"1100011001111" WHEN "0010000100",
"0100001101010" WHEN "0010000101",
"0011001010101" WHEN "0010000110",
"0101111001001" WHEN "0010000111",
"0010100110111" WHEN "0010001000",
"1001001101111" WHEN "0010001001",
"1101101000100" WHEN "0010001010",
"1010000101011" WHEN "0010001011",
"0001110100110" WHEN "0010001100",
"0000000001111" WHEN "0010001101",
"0001001100001" WHEN "0010001110",
"0111000110010" WHEN "0010001111",
"0100100000100" WHEN "0010010000",
"0000111101011" WHEN "0010010001",
"1100000011101" WHEN "0010010010",
"1101010010110" WHEN "0010010011",
"1011010100111" WHEN "0010010100",
"1110110100010" WHEN "0010010101",
"0010000011000" WHEN "0010010110",
"0101001101100" WHEN "0010010111",
"1100101000100" WHEN "0010011000",
"1000100010110" WHEN "0010011001",
"1111000110100" WHEN "0010011010",
"0011001101100" WHEN "0010011011",
"0111001111111" WHEN "0010011100",
"1001010011110" WHEN "0010011101",
"0001000101001" WHEN "0010011110",
"0010110111000" WHEN "0010011111",
"0111010011001" WHEN "0010100000",
"1111010111011" WHEN "0010100001",
"0001001101010" WHEN "0010100010",
"0000010100101" WHEN "0010100011",
"1000001110111" WHEN "0010100100",
"1100000001100" WHEN "0010100101",
"0110010011001" WHEN "0010100110",
"1110011100010" WHEN "0010100111",
"1000010001101" WHEN "0010101000",
"1001110101011" WHEN "0010101001",
"1110001011000" WHEN "0010101010",
"1001000010111" WHEN "0010101011",
"0111000001111" WHEN "0010101100",
"0001000110101" WHEN "0010101101",
"0110011010000" WHEN "0010101110",
"1100011000101" WHEN "0010101111",
"1010111011110" WHEN "0010110000",
"1110100111100" WHEN "0010110001",
"1010111001110" WHEN "0010110010",
"1100100110101" WHEN "0010110011",
"0111111000101" WHEN "0010110100",
"1100011110111" WHEN "0010110101",
"0011011010100" WHEN "0010110110",
"0010010111110" WHEN "0010110111",
"1100010000000" WHEN "0010111000",
"1001101111001" WHEN "0010111001",
"0000100010101" WHEN "0010111010",
"0100110111100" WHEN "0010111011",
"0001000100011" WHEN "0010111100",
"1010011010111" WHEN "0010111101",
"0100011010010" WHEN "0010111110",
"0100100100001" WHEN "0010111111",
"1110010000001" WHEN "0011000000",
"0111100011010" WHEN "0011000001",
"0011100001100" WHEN "0011000010",
"1110001110100" WHEN "0011000011",
"0100000110000" WHEN "0011000100",
"0100011101100" WHEN "0011000101",
"1111000011111" WHEN "0011000110",
"1001111010000" WHEN "0011000111",
"1000011010110" WHEN "0011001000",
"1101101101111" WHEN "0011001001",
"0011001001011" WHEN "0011001010",
"1110100101001" WHEN "0011001011",
"1111001110001" WHEN "0011001100",
"0100111001001" WHEN "0011001101",
"0001011000011" WHEN "0011001110",
"0000100011010" WHEN "0011001111",
"1100101010010" WHEN "0011010000",
"1100001010001" WHEN "0011010001",
"0010001100100" WHEN "0011010010",
"0110011110110" WHEN "0011010011",
"0000110010010" WHEN "0011010100",
"0100110000100" WHEN "0011010101",
"1110010110110" WHEN "0011010110",
"1111011111101" WHEN "0011010111",
"1100011000111" WHEN "0011011000",
"0100001000010" WHEN "0011011001",
"1101001100110" WHEN "0011011010",
"1011100000101" WHEN "0011011011",
"1001111010000" WHEN "0011011100",
"0100011110111" WHEN "0011011101",
"0011111110010" WHEN "0011011110",
"0110011101110" WHEN "0011011111",
"1101010001000" WHEN "0011100000",
"0111011011010" WHEN "0011100001",
"0110110111111" WHEN "0011100010",
"1110111100101" WHEN "0011100011",
"0010001010011" WHEN "0011100100",
"0011001100000" WHEN "0011100101",
"0101001101100" WHEN "0011100110",
"0001000111111" WHEN "0011100111",
"0001001011110" WHEN "0011101000",
"0101110100010" WHEN "0011101001",
"0111010011101" WHEN "0011101010",
"0111110010001" WHEN "0011101011",
"0001110001111" WHEN "0011101100",
"1100101111001" WHEN "0011101101",
"0110100101000" WHEN "0011101110",
"0110101010100" WHEN "0011101111",
"1001000011100" WHEN "0011110000",
"0010101111000" WHEN "0011110001",
"1110011110011" WHEN "0011110010",
"1011001010001" WHEN "0011110011",
"1011111001011" WHEN "0011110100",
"1010100110110" WHEN "0011110101",
"1111101110110" WHEN "0011110110",
"0010110110011" WHEN "0011110111",
"1101111100111" WHEN "0011111000",
"0001010011111" WHEN "0011111001",
"1110100111111" WHEN "0011111010",
"0010010001001" WHEN "0011111011",
"0110011110101" WHEN "0011111100",
"0111100110101" WHEN "0011111101",
"1000110000011" WHEN "0011111110",
"1001100100001" WHEN "0011111111",
"0000000000000" when others;
end behavioural;
