--Splits a 7 bit binary signal into 2
--BCD coded signals
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity Bit7ToBCD is
    port( BIn : in STD_LOGIC_VECTOR( 6 downto 0 );
           MSD, LSD: out STD_LOGIC_VECTOR( 3 downto 0 ));
end Bit7ToBCD;

architecture behavioural of Bit7ToBCD is

begin
    --Generated with BCDgen.java 
	with BIn select
	MSD <= "0000" WHEN "0000000",
			"0000" WHEN "0000001",
			"0000" WHEN "0000010",
			"0000" WHEN "0000011",
			"0000" WHEN "0000100",
			"0000" WHEN "0000101",
			"0000" WHEN "0000110",
			"0000" WHEN "0000111",
			"0000" WHEN "0001000",
			"0000" WHEN "0001001",
			"0001" WHEN "0001010",
			"0001" WHEN "0001011",
			"0001" WHEN "0001100",
			"0001" WHEN "0001101",
			"0001" WHEN "0001110",
			"0001" WHEN "0001111",
			"0001" WHEN "0010000",
			"0001" WHEN "0010001",
			"0001" WHEN "0010010",
			"0001" WHEN "0010011",
			"0010" WHEN "0010100",
			"0010" WHEN "0010101",
			"0010" WHEN "0010110",
			"0010" WHEN "0010111",
			"0010" WHEN "0011000",
			"0010" WHEN "0011001",
			"0010" WHEN "0011010",
			"0010" WHEN "0011011",
			"0010" WHEN "0011100",
			"0010" WHEN "0011101",
			"0011" WHEN "0011110",
			"0011" WHEN "0011111",
			"0011" WHEN "0100000",
			"0011" WHEN "0100001",
			"0011" WHEN "0100010",
			"0011" WHEN "0100011",
			"0011" WHEN "0100100",
			"0011" WHEN "0100101",
			"0011" WHEN "0100110",
			"0011" WHEN "0100111",
			"0100" WHEN "0101000",
			"0100" WHEN "0101001",
			"0100" WHEN "0101010",
			"0100" WHEN "0101011",
			"0100" WHEN "0101100",
			"0100" WHEN "0101101",
			"0100" WHEN "0101110",
			"0100" WHEN "0101111",
			"0100" WHEN "0110000",
			"0100" WHEN "0110001",
			"0101" WHEN "0110010",
			"0101" WHEN "0110011",
			"0101" WHEN "0110100",
			"0101" WHEN "0110101",
			"0101" WHEN "0110110",
			"0101" WHEN "0110111",
			"0101" WHEN "0111000",
			"0101" WHEN "0111001",
			"0101" WHEN "0111010",
			"0101" WHEN "0111011",
			"0110" WHEN "0111100",
			"0110" WHEN "0111101",
			"0110" WHEN "0111110",
			"0110" WHEN "0111111",
			"0110" WHEN "1000000",
			"0110" WHEN "1000001",
			"0110" WHEN "1000010",
			"0110" WHEN "1000011",
			"0110" WHEN "1000100",
			"0110" WHEN "1000101",
			"0111" WHEN "1000110",
			"0111" WHEN "1000111",
			"0111" WHEN "1001000",
			"0111" WHEN "1001001",
			"0111" WHEN "1001010",
			"0111" WHEN "1001011",
			"0111" WHEN "1001100",
			"0111" WHEN "1001101",
			"0111" WHEN "1001110",
			"0111" WHEN "1001111",
			"1000" WHEN "1010000",
			"1000" WHEN "1010001",
			"1000" WHEN "1010010",
			"1000" WHEN "1010011",
			"1000" WHEN "1010100",
			"1000" WHEN "1010101",
			"1000" WHEN "1010110",
			"1000" WHEN "1010111",
			"1000" WHEN "1011000",
			"1000" WHEN "1011001",
			"1001" WHEN "1011010",
			"1001" WHEN "1011011",
			"1001" WHEN "1011100",
			"1001" WHEN "1011101",
			"1001" WHEN "1011110",
			"1001" WHEN "1011111",
			"1001" WHEN "1100000",
			"1001" WHEN "1100001",
			"1001" WHEN "1100010",
			"1001" WHEN "1100011",
			"1111" WHEN OTHERS;
	with BIn select
	LSD <= "0000" WHEN "0000000",
				"0001" WHEN "0000001",
				"0010" WHEN "0000010",
				"0011" WHEN "0000011",
				"0100" WHEN "0000100",
				"0101" WHEN "0000101",
				"0110" WHEN "0000110",
				"0111" WHEN "0000111",
				"1000" WHEN "0001000",
				"1001" WHEN "0001001",
				"0000" WHEN "0001010",
				"0001" WHEN "0001011",
				"0010" WHEN "0001100",
				"0011" WHEN "0001101",
				"0100" WHEN "0001110",
				"0101" WHEN "0001111",
				"0110" WHEN "0010000",
				"0111" WHEN "0010001",
				"1000" WHEN "0010010",
				"1001" WHEN "0010011",
				"0000" WHEN "0010100",
				"0001" WHEN "0010101",
				"0010" WHEN "0010110",
				"0011" WHEN "0010111",
				"0100" WHEN "0011000",
				"0101" WHEN "0011001",
				"0110" WHEN "0011010",
				"0111" WHEN "0011011",
				"1000" WHEN "0011100",
				"1001" WHEN "0011101",
				"0000" WHEN "0011110",
				"0001" WHEN "0011111",
				"0010" WHEN "0100000",
				"0011" WHEN "0100001",
				"0100" WHEN "0100010",
				"0101" WHEN "0100011",
				"0110" WHEN "0100100",
				"0111" WHEN "0100101",
				"1000" WHEN "0100110",
				"1001" WHEN "0100111",
				"0000" WHEN "0101000",
				"0001" WHEN "0101001",
				"0010" WHEN "0101010",
				"0011" WHEN "0101011",
				"0100" WHEN "0101100",
				"0101" WHEN "0101101",
				"0110" WHEN "0101110",
				"0111" WHEN "0101111",
				"1000" WHEN "0110000",
				"1001" WHEN "0110001",
				"0000" WHEN "0110010",
				"0001" WHEN "0110011",
				"0010" WHEN "0110100",
				"0011" WHEN "0110101",
				"0100" WHEN "0110110",
				"0101" WHEN "0110111",
				"0110" WHEN "0111000",
				"0111" WHEN "0111001",
				"1000" WHEN "0111010",
				"1001" WHEN "0111011",
				"0000" WHEN "0111100",
				"0001" WHEN "0111101",
				"0010" WHEN "0111110",
				"0011" WHEN "0111111",
				"0100" WHEN "1000000",
				"0101" WHEN "1000001",
				"0110" WHEN "1000010",
				"0111" WHEN "1000011",
				"1000" WHEN "1000100",
				"1001" WHEN "1000101",
				"0000" WHEN "1000110",
				"0001" WHEN "1000111",
				"0010" WHEN "1001000",
				"0011" WHEN "1001001",
				"0100" WHEN "1001010",
				"0101" WHEN "1001011",
				"0110" WHEN "1001100",
				"0111" WHEN "1001101",
				"1000" WHEN "1001110",
				"1001" WHEN "1001111",
				"0000" WHEN "1010000",
				"0001" WHEN "1010001",
				"0010" WHEN "1010010",
				"0011" WHEN "1010011",
				"0100" WHEN "1010100",
				"0101" WHEN "1010101",
				"0110" WHEN "1010110",
				"0111" WHEN "1010111",
				"1000" WHEN "1011000",
				"1001" WHEN "1011001",
				"0000" WHEN "1011010",
				"0001" WHEN "1011011",
				"0010" WHEN "1011100",
				"0011" WHEN "1011101",
				"0100" WHEN "1011110",
				"0101" WHEN "1011111",
				"0110" WHEN "1100000",
				"0111" WHEN "1100001",
				"1000" WHEN "1100010",
				"1001" WHEN "1100011",
				"1111" WHEN OTHERS;
	
end behavioural;
    
