library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity diet_rom is
    port(   addr : in std_logic_vector( 6 downto 0 );
            do : out std_logic_vector( 3 downto 0 ) );
end diet_rom;

architecture behavioural of diet_rom is
begin
    with addr select
    do <= "0000" WHEN "0000000",
            "0000" WHEN "0000001",
            "0000" WHEN "0000010",
            "0000" WHEN "0000011",
            "0000" WHEN "0000100",
            "0000" WHEN "0000101",
            "0000" WHEN "0000110",
            "0000" WHEN "0000111",
            "0000" WHEN "0001000",
            "0000" WHEN "0001001",
            "0001" WHEN "0001010",
            "0001" WHEN "0001011",
            "0001" WHEN "0001100",
            "0001" WHEN "0001101",
            "0001" WHEN "0001110",
            "0001" WHEN "0001111",
            "0001" WHEN "0010000",
            "0001" WHEN "0010001",
            "0001" WHEN "0010010",
            "0001" WHEN "0010011",
            "0010" WHEN "0010100",
            "0010" WHEN "0010101",
            "0010" WHEN "0010110",
            "0010" WHEN "0010111",
            "0010" WHEN "0011000",
            "0010" WHEN "0011001",
            "0010" WHEN "0011010",
            "0010" WHEN "0011011",
            "0010" WHEN "0011100",
            "0010" WHEN "0011101",
            "0011" WHEN "0011110",
            "0011" WHEN "0011111",
            "0011" WHEN "0100000",
            "0011" WHEN "0100001",
            "0011" WHEN "0100010",
            "0011" WHEN "0100011",
            "0011" WHEN "0100100",
            "0011" WHEN "0100101",
            "0011" WHEN "0100110",
            "0011" WHEN "0100111",
            "0100" WHEN "0101000",
            "0100" WHEN "0101001",
            "0100" WHEN "0101010",
            "0100" WHEN "0101011",
            "0100" WHEN "0101100",
            "0100" WHEN "0101101",
            "0100" WHEN "0101110",
            "0100" WHEN "0101111",
            "0100" WHEN "0110000",
            "0100" WHEN "0110001",
            "0101" WHEN "0110010",
            "0101" WHEN "0110011",
            "0101" WHEN "0110100",
            "0101" WHEN "0110101",
            "0101" WHEN "0110110",
            "0101" WHEN "0110111",
            "0101" WHEN "0111000",
            "0101" WHEN "0111001",
            "0101" WHEN "0111010",
            "0101" WHEN "0111011",
            "0110" WHEN "0111100",
            "0110" WHEN "0111101",
            "0110" WHEN "0111110",
            "0110" WHEN "0111111",
            "0110" WHEN "1000000",
            "0110" WHEN "1000001",
            "0110" WHEN "1000010",
            "0110" WHEN "1000011",
            "0110" WHEN "1000100",
            "0110" WHEN "1000101",
            "0111" WHEN "1000110",
            "0111" WHEN "1000111",
            "0111" WHEN "1001000",
            "0111" WHEN "1001001",
            "0111" WHEN "1001010",
            "0111" WHEN "1001011",
            "0111" WHEN "1001100",
            "0111" WHEN "1001101",
            "0111" WHEN "1001110",
            "0111" WHEN "1001111",
            "1000" WHEN "1010000",
            "1000" WHEN "1010001",
            "1000" WHEN "1010010",
            "1000" WHEN "1010011",
            "1000" WHEN "1010100",
            "1000" WHEN "1010101",
            "1000" WHEN "1010110",
            "1000" WHEN "1010111",
            "1000" WHEN "1011000",
            "1000" WHEN "1011001",
            "1001" WHEN "1011010",
            "1001" WHEN "1011011",
            "1001" WHEN "1011100",
            "1001" WHEN "1011101",
            "1001" WHEN "1011110",
            "1001" WHEN "1011111",
            "1001" WHEN "1100000",
            "1001" WHEN "1100001",
            "1001" WHEN "1100010",
            "1001" WHEN "1100011",
            "1111" WHEN OTHERS;
end behavioural;

