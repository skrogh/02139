library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity diet_rom is
    port(   addr : in std_logic_vector( 7 downto 0 );
            do : out std_logic_vector( 7 downto 0 ) );
end diet_rom;

architecture behavioural of diet_rom is
begin
    with addr select
    do <= "11000110" WHEN "00000000",
"01000100" WHEN "00000001",
"01010111" WHEN "00000010",
"10100011" WHEN "00000011",
"01101001" WHEN "00000100",
"01100000" WHEN "00000101",
"10000101" WHEN "00000110",
"11101100" WHEN "00000111",
"01001001" WHEN "00001000",
"11100010" WHEN "00001001",
"11010001" WHEN "00001010",
"00010010" WHEN "00001011",
"01110110" WHEN "00001100",
"11000011" WHEN "00001101",
"00011000" WHEN "00001110",
"01000011" WHEN "00001111",
"11111010" WHEN "00010000",
"11001000" WHEN "00010001",
"11000000" WHEN "00010010",
"11010100" WHEN "00010011",
"10000110" WHEN "00010100",
"01111101" WHEN "00010101",
"11000001" WHEN "00010110",
"01101111" WHEN "00010111",
"01000000" WHEN "00011000",
"10110010" WHEN "00011001",
"01100010" WHEN "00011010",
"01111010" WHEN "00011011",
"11101001" WHEN "00011100",
"10101101" WHEN "00011101",
"00010001" WHEN "00011110",
"00001010" WHEN "00011111",
"01101000" WHEN "00100000",
"01101010" WHEN "00100001",
"00010010" WHEN "00100010",
"01101000" WHEN "00100011",
"11001010" WHEN "00100100",
"00010111" WHEN "00100101",
"11101011" WHEN "00100110",
"01001111" WHEN "00100111",
"10000010" WHEN "00101000",
"01000011" WHEN "00101001",
"10011011" WHEN "00101010",
"00000101" WHEN "00101011",
"01110101" WHEN "00101100",
"01111101" WHEN "00101101",
"11000010" WHEN "00101110",
"11011110" WHEN "00101111",
"11101111" WHEN "00110000",
"10111000" WHEN "00110001",
"10101101" WHEN "00110010",
"00010010" WHEN "00110011",
"00110101" WHEN "00110100",
"01001100" WHEN "00110101",
"00111111" WHEN "00110110",
"10000010" WHEN "00110111",
"10111011" WHEN "00111000",
"01101000" WHEN "00111001",
"01001011" WHEN "00111010",
"10110010" WHEN "00111011",
"01111011" WHEN "00111100",
"10010001" WHEN "00111101",
"10111010" WHEN "00111110",
"01000000" WHEN "00111111",
"00000101" WHEN "01000000",
"00010110" WHEN "01000001",
"01001110" WHEN "01000010",
"00100010" WHEN "01000011",
"00101011" WHEN "01000100",
"01111000" WHEN "01000101",
"01100010" WHEN "01000110",
"00111011" WHEN "01000111",
"00000111" WHEN "01001000",
"01111000" WHEN "01001001",
"01100000" WHEN "01001010",
"00110111" WHEN "01001011",
"01001111" WHEN "01001100",
"10110110" WHEN "01001101",
"11101110" WHEN "01001110",
"00100111" WHEN "01001111",
"10000101" WHEN "01010000",
"11110100" WHEN "01010001",
"00000011" WHEN "01010010",
"00001011" WHEN "01010011",
"10001110" WHEN "01010100",
"10011111" WHEN "01010101",
"00110101" WHEN "01010110",
"01010111" WHEN "01010111",
"10111110" WHEN "01011000",
"10001101" WHEN "01011001",
"10001010" WHEN "01011010",
"01111100" WHEN "01011011",
"00100000" WHEN "01011100",
"11100100" WHEN "01011101",
"00001100" WHEN "01011110",
"10101100" WHEN "01011111",
"00011001" WHEN "01100000",
"10110011" WHEN "01100001",
"00011001" WHEN "01100010",
"01101001" WHEN "01100011",
"00011100" WHEN "01100100",
"00011000" WHEN "01100101",
"01000001" WHEN "01100110",
"11100011" WHEN "01100111",
"00101001" WHEN "01101000",
"10101001" WHEN "01101001",
"00001101" WHEN "01101010",
"11001010" WHEN "01101011",
"01100101" WHEN "01101100",
"10001000" WHEN "01101101",
"10011100" WHEN "01101110",
"00010001" WHEN "01101111",
"11010001" WHEN "01110000",
"10110011" WHEN "01110001",
"01110001" WHEN "01110010",
"00000110" WHEN "01110011",
"10001010" WHEN "01110100",
"00010000" WHEN "01110101",
"00110011" WHEN "01110110",
"01000100" WHEN "01110111",
"10010100" WHEN "01111000",
"01001111" WHEN "01111001",
"01001000" WHEN "01111010",
"00111110" WHEN "01111011",
"01010110" WHEN "01111100",
"11011011" WHEN "01111101",
"01111101" WHEN "01111110",
"10100100" WHEN "01111111",
"01011101" WHEN "10000000",
"00010001" WHEN "10000001",
"11011101" WHEN "10000010",
"01010110" WHEN "10000011",
"11110100" WHEN "10000100",
"01011000" WHEN "10000101",
"11110011" WHEN "10000110",
"01111001" WHEN "10000111",
"01001111" WHEN "10001000",
"00000101" WHEN "10001001",
"01110011" WHEN "10001010",
"11111010" WHEN "10001011",
"11100000" WHEN "10001100",
"11000000" WHEN "10001101",
"00110000" WHEN "10001110",
"00000010" WHEN "10001111",
"01101001" WHEN "10010000",
"10010000" WHEN "10010001",
"11100000" WHEN "10010010",
"11110110" WHEN "10010011",
"00000000" WHEN "10010100",
"11111000" WHEN "10010101",
"11001101" WHEN "10010110",
"11111011" WHEN "10010111",
"00001001" WHEN "10011000",
"01000110" WHEN "10011001",
"00010001" WHEN "10011010",
"10001010" WHEN "10011011",
"10100100" WHEN "10011100",
"10110110" WHEN "10011101",
"01111111" WHEN "10011110",
"00110100" WHEN "10011111",
"10100000" WHEN "10100000",
"00101111" WHEN "10100001",
"01101110" WHEN "10100010",
"10100001" WHEN "10100011",
"01010010" WHEN "10100100",
"00011101" WHEN "10100101",
"00101011" WHEN "10100110",
"10110110" WHEN "10100111",
"00011100" WHEN "10101000",
"01011110" WHEN "10101001",
"10011011" WHEN "10101010",
"00001111" WHEN "10101011",
"01111111" WHEN "10101100",
"01010101" WHEN "10101101",
"11110011" WHEN "10101110",
"00101011" WHEN "10101111",
"11011001" WHEN "10110000",
"11101110" WHEN "10110001",
"00011110" WHEN "10110010",
"00101111" WHEN "10110011",
"11000010" WHEN "10110100",
"11000011" WHEN "10110101",
"01101111" WHEN "10110110",
"10101010" WHEN "10110111",
"00110001" WHEN "10111000",
"10110011" WHEN "10111001",
"11010110" WHEN "10111010",
"10100101" WHEN "10111011",
"00001010" WHEN "10111100",
"11011000" WHEN "10111101",
"10100011" WHEN "10111110",
"00010110" WHEN "10111111",
"11011101" WHEN "11000000",
"00111110" WHEN "11000001",
"01010000" WHEN "11000010",
"11111111" WHEN "11000011",
"11011000" WHEN "11000100",
"10111100" WHEN "11000101",
"01010101" WHEN "11000110",
"10011100" WHEN "11000111",
"11010110" WHEN "11001000",
"11111111" WHEN "11001001",
"01101001" WHEN "11001010",
"10000011" WHEN "11001011",
"10101100" WHEN "11001100",
"00110010" WHEN "11001101",
"11010111" WHEN "11001110",
"00011010" WHEN "11001111",
"01100000" WHEN "11010000",
"10100010" WHEN "11010001",
"11001001" WHEN "11010010",
"01101101" WHEN "11010011",
"00000101" WHEN "11010100",
"01111100" WHEN "11010101",
"01110011" WHEN "11010110",
"01101010" WHEN "11010111",
"01101110" WHEN "11011000",
"11110100" WHEN "11011001",
"00100010" WHEN "11011010",
"01011011" WHEN "11011011",
"10101100" WHEN "11011100",
"00110001" WHEN "11011101",
"11111110" WHEN "11011110",
"11100001" WHEN "11011111",
"10010010" WHEN "11100000",
"11110011" WHEN "11100001",
"01000100" WHEN "11100010",
"10111110" WHEN "11100011",
"00101111" WHEN "11100100",
"00110000" WHEN "11100101",
"01001011" WHEN "11100110",
"01111101" WHEN "11100111",
"00010000" WHEN "11101000",
"11001010" WHEN "11101001",
"01110001" WHEN "11101010",
"01110110" WHEN "11101011",
"11000101" WHEN "11101100",
"00110001" WHEN "11101101",
"01111100" WHEN "11101110",
"10001110" WHEN "11101111",
"11100010" WHEN "11110000",
"11011111" WHEN "11110001",
"01111001" WHEN "11110010",
"00001010" WHEN "11110011",
"11110110" WHEN "11110100",
"10100110" WHEN "11110101",
"01110001" WHEN "11110110",
"11011001" WHEN "11110111",
"10111101" WHEN "11111000",
"01000001" WHEN "11111001",
"10011001" WHEN "11111010",
"00001100" WHEN "11111011",
"11000110" WHEN "11111100",
"11011001" WHEN "11111101",
"11001011" WHEN "11111110",
"10000100" WHEN "11111111",
            "11111111" WHEN OTHERS;
end behavioural;

