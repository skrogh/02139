library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
entity rom is
port( addr : in std_logic_vector( 9 downto 0 );
do : out std_logic_vector( 12 downto 0 ) );
end rom;
architecture behavioural of rom is
begin
with addr select
do <= "0111011111111" WHEN "0000000000",
"0110110100000" WHEN "0000000001",
"0111100000000" WHEN "0000000010",
"1000100000001" WHEN "0000000011",
"0111100000001" WHEN "0000000100",
"1000100000010" WHEN "0000000101",
"0111100000010" WHEN "0000000110",
"1000100000100" WHEN "0000000111",
"0111100000011" WHEN "0000001000",
"1000100001000" WHEN "0000001001",
"0111100000100" WHEN "0000001010",
"1000100010000" WHEN "0000001011",
"0111100000101" WHEN "0000001100",
"1000100100000" WHEN "0000001101",
"0111100000110" WHEN "0000001110",
"1000101000000" WHEN "0000001111",
"0111100000111" WHEN "0000010000",
"1000110000000" WHEN "0000010001",
"0111100001000" WHEN "0000010010",
"1000111110000" WHEN "0000010011",
"0111100001001" WHEN "0000010100",
"1000100001111" WHEN "0000010101",
"0010101000000" WHEN "0000010110",
"0111000000001" WHEN "0000010111",
"0011000010000" WHEN "0000011000",
"0010100110000" WHEN "0000011001",
"0010100100000" WHEN "0000011010",
"0000100100001" WHEN "0000011011",
"0101000000010" WHEN "0000011100",
"0100100000010" WHEN "0000011101",
"0000100110001" WHEN "0000011110",
"0101000000010" WHEN "0000011111",
"0100100000110" WHEN "0000100000",
"1000001000000" WHEN "0000100001",
"0000101000001" WHEN "0000100010",
"1001101010000" WHEN "0000100011",
"0110110100101" WHEN "0000100100",
"0110001010001" WHEN "0000100101",
"0111000000001" WHEN "0000100110",
"1010001010000" WHEN "0000100111",
"0001001010001" WHEN "0000101000",
"0101000000010" WHEN "0000101001",
"0100100000101" WHEN "0000101010",
"0110001010001" WHEN "0000101011",
"0111000000001" WHEN "0000101100",
"1010001010000" WHEN "0000101101",
"0001001010001" WHEN "0000101110",
"0101100000100" WHEN "0000101111",
"0100100010010" WHEN "0000110000",
"0000000000000" when others;
end behavioural;
