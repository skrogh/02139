library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
entity rom is
port( clk : in std_logic;
addr : in std_logic_vector( 9 downto 0 );
do : out std_logic_vector( 12 downto 0 ) );
end rom;
architecture behavioural of rom is
signal addr_clkd : std_logic_vector( 9 downto 0 );
begin
process( CLK ) begin
if rising_edge( CLK ) then
addr_clkd <= addr;
end if;
end process;
with addr_clkd select
do <= "0000000000000" WHEN "0000000000",
"0111001001111" WHEN "0000000001",
"0010000010110" WHEN "0000000010",
"0001100010100" WHEN "0000000011",
"0011000100000" WHEN "0000000100",
"1010100000001" WHEN "0000000101",
"0000100000001" WHEN "0000000110",
"1010100000001" WHEN "0000000111",
"0001000000001" WHEN "0000001000",
"0010100000000" WHEN "0000001001",
"0001000000001" WHEN "0000001010",
"0000000000000" WHEN "0000001011",
"0011100001110" WHEN "0000001100",
"0100000000010" WHEN "0000001101",
"0100100000001" WHEN "0000001110",
"0000000000000" WHEN "0000001111",
"1011100110000" WHEN "0000010000",
"1100001000000" WHEN "0000010001",
"0111000000001" WHEN "0000010010",
"0000100110000" WHEN "0000010011",
"0111000001000" WHEN "0000010100",
"0000100110000" WHEN "0000010101",
"0010100000000" WHEN "0000010110",
"1010101000000" WHEN "0000010111",
"0100000000011" WHEN "0000011000",
"0111011111111" WHEN "0000011001",
"0100100000001" WHEN "0000011010",
"0111000000001" WHEN "0000011011",
"0011000010000" WHEN "0000011100",
"1011000010000" WHEN "0000011101",
"0101011111111" WHEN "0000011110",
"1011000000000" WHEN "0000011111",
"0101111111111" WHEN "0000100000",
"1011000000001" WHEN "0000100001",
"0101000000101" WHEN "0000100010",
"0000000000000" WHEN "0000100011",
"0000000000000" WHEN "0000100100",
"0000000000000" WHEN "0000100101",
"0100000000010" WHEN "0000100110",
"0101100000001" WHEN "0000100111",
"0111011111111" WHEN "0000101000",
"0110100000000" WHEN "0000101001",
"0110101110000" WHEN "0000101010",
"0010100000000" WHEN "0000101011",
"0110000000111" WHEN "0000101100",
"0110000000000" WHEN "0000101101",
"0111100000001" WHEN "0000101110",
"1000111110000" WHEN "0000101111",
"0111000001111" WHEN "0000110000",
"1001000000000" WHEN "0000110001",
"0111000000010" WHEN "0000110010",
"1000000000000" WHEN "0000110011",
"1001000000000" WHEN "0000110100",
"1001100010000" WHEN "0000110101",
"1100101000011" WHEN "0000110110",
"0000000000000" when others;
end behavioural;
